`ifndef __SSW_INFO_H__
`define __SSW_INFO_H__


`define STACK_SIZE (32'h 2000)
`define DATA_ALIGN_SIZE 4
`define PRINTF_USING_UART
//`define PRINTF_USING_OLED
`define TEMPORARY_CACHING_HEAP_START 0
`define TEMPORARY_CACHING_HEAP_SIZE 0
`define TEMPORARY_CACHING_HEAP_LAST 0
`define NUM_THREAD_PER_TEAM 1
`define UNCACHEABLE_MEMORY_REGION sram
`define CACHEABLE_MEMORY_REGION sram
`define BIGDATA_MEMORY_REGION sram

`endif