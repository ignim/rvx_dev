/*****************/
/* Custom Region */
/*****************/

// wire spi_common_sclk;
// wire spi_common_sdq0;
// wire clk_system;
// wire clk_core;
// wire clk_system_external;
// wire clk_system_debug;
// wire clk_local_access;
// wire clk_process_000;
// wire clk_noc;
// wire clk_sdram_cell;
// wire clk_sdram_if;
// wire gclk_system;
// wire gclk_core;
// wire gclk_system_external;
// wire gclk_system_debug;
// wire gclk_local_access;
// wire gclk_process_000;
// wire gclk_noc;
// wire gclk_sdram_cell;
// wire gclk_sdram_if;
// wire tick_1us;
// wire tick_62d5ms;
// wire tick_gpio;
// wire global_rstnn;
// wire global_rstpp;
// wire [(6)-1:0] rstnn_seqeunce;
// wire [(6)-1:0] rstpp_seqeunce;
// wire rstnn_user;
// wire rstpp_user;

/* DO NOT MODIFY THE ABOVE */
/* MUST MODIFY THE BELOW   */
