`ifndef __HW_INFO_H__
`define __HW_INFO_H__


`define NUM_CORE_USER 1
`define NUM_CORE_TEAM 1
`define NUM_LOCK_USER 0
`define NUM_LOCK_SYSTEM 0
`define NUM_BARRIER_USER 0
`define NUM_BARRIER_SYSTEM 0
`define NUM_AUTO_ID 0
`define NUM_GLOBAL_TAG 0
`define SRAM_SIZE (32'h 20000)
`define SRAM_CELL_SIZE (32'h 20000)
`define DRAM_SIZE 0
`define INCLUDE_IROM
`define SYSTEM_CLK_HZ 50000000
`define CORE_CLK_HZ 50000000
`define UART_CLK_HZ 50000000
`define SPI_CLK_HZ 50000000
`define I2C_CLK_HZ 50000000
`define OLED_CLK_HZ 50000000
`define TICK_HZ 1000000
`define NUM_UART_READYMADE 1
`define NUM_SPI_READYMADE 1
`define NUM_I2C_READYMADE 1
`define NUM_GPIO_READYMADE 0
`define NUM_UART_USER 0
`define NUM_SPI_USER 0
`define NUM_I2C_USER 0
`define NUM_GPIO_USER 0
`define NUM_LED_CHECKER 1
`define NUM_AIOIF 0
`define NUM_SWITCH_SLIDE_READYMADE 0
`define INCLUDE_SRAM
//`define INCLUDE_SLOW_DRAM
//`define INCLUDE_FAST_DRAM
//`define INCLUDE_DRAM
`define INCLUDE_BOOT_MODE
//`define INCLUDE_CACHE
`define INCLUDE_TIMER
//`define INCLUDE_PLIC
//`define INCLUDE_CORE_JTAG
`define INCLUDE_OLED
`define INCLUDE_OLED_BW
`define INCLUDE_OLED_RGB
`define INCLUDE_SPI_FLASH
//`define INCLUDE_VIDEO
`define INCLUDE_UART_PRINTF
//`define INCLUDE_OLEDBW_PRINTF
//`define INCLUDE_FUSE_BOX
//`define INCLUDE_USER_INTERRUPTS
//`define INCLUDE_ARDUCAM
//`define INCLUDE_BLUETOOTH
//`define INCLUDE_WIFI
//`define INCLUDE_JPEG_ENCODER
//`define INCLUDE_JPEGLS_ENCODER
//`define INCLUDE_HBC1_TX
//`define INCLUDE_HBC1_RX
`define INCLUDE_CORE_PERI_GROUP
//`define USE_NOC_DEBUG
//`define USE_TEMPORARY_CACHING
//`define USE_SW_BARRIER
`define USE_HW_BARRIER
`define USE_PROFILING
`define NOC_FLIT_DIVISOR 1
`define PLATFORM_NAME "tip_arty"
`define INCLUDE_RVC_ORCA
`define NUM_CORE 1
`define NUM_REAL_CORE 1
//`define USE_MULTICORE
`define NUM_BARRIER 0
`define NUM_LOCK 0
`define SPI_INDEX_FOR_READYMADE 0
`define SPI_INDEX_FOR_USER 1
`define SPI_INDEX_FOR_SYSTEM 1
`define SPI_INDEX_FOR_AIOIF 1
`define SPI_INDEX_FOR_OLED 1
`define SPI_INDEX_FOR_SPI_FLASH 2
`define NUM_SPI_SYSTEM 2
`define UART_INDEX_FOR_READYMADE 0
`define UART_INDEX_FOR_USER 1
`define UART_INDEX_FOR_SYSTEM 1
`define UART_INDEX_FOR_AIOIF 1
`define UART_INDEX_FOR_UART_PRINTF 1
`define NUM_UART_SYSTEM 1
`define I2C_INDEX_FOR_READYMADE 0
`define I2C_INDEX_FOR_USER 1
`define I2C_INDEX_FOR_SYSTEM 1
`define I2C_INDEX_FOR_AIOIF 1
`define NUM_I2C_SYSTEM 0
`define GPIO_INDEX_FOR_READYMADE 0
`define GPIO_INDEX_FOR_USER 0
`define GPIO_INDEX_FOR_SYSTEM 0
`define GPIO_INDEX_FOR_AIOIF 0
`define GPIO_INDEX_FOR_SWITCH_SLIDE_READYMADE 0
`define NUM_GPIO_SYSTEM 0
`define SRAM_ADDR (32'h 40000000)
`define APP_ADDR (32'h 40000000)
`define NUM_UART 2
`define NUM_SPI 3
`define NUM_I2C 1
`define NUM_GPIO 0
`define INCLUDE_CORE_USER
`define INCLUDE_CORE_TEAM
//`define INCLUDE_LOCK_USER
//`define INCLUDE_LOCK_SYSTEM
//`define INCLUDE_BARRIER_USER
//`define INCLUDE_BARRIER_SYSTEM
//`define INCLUDE_AUTO_ID
//`define INCLUDE_GLOBAL_TAG
`define INCLUDE_UART_READYMADE
`define INCLUDE_SPI_READYMADE
`define INCLUDE_I2C_READYMADE
//`define INCLUDE_GPIO_READYMADE
//`define INCLUDE_UART_USER
//`define INCLUDE_SPI_USER
//`define INCLUDE_I2C_USER
//`define INCLUDE_GPIO_USER
`define INCLUDE_LED_CHECKER
//`define INCLUDE_AIOIF
//`define INCLUDE_SWITCH_SLIDE_READYMADE
`define INCLUDE_CORE
`define INCLUDE_REAL_CORE
//`define INCLUDE_BARRIER
//`define INCLUDE_LOCK
`define INCLUDE_SPI_SYSTEM
`define INCLUDE_UART_SYSTEM
//`define INCLUDE_I2C_SYSTEM
//`define INCLUDE_GPIO_SYSTEM
`define INCLUDE_UART
`define INCLUDE_SPI
`define INCLUDE_I2C
//`define INCLUDE_GPIO
`define NUM_PREDEFINED_CLOCK 0

`endif