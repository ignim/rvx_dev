`ifndef __MEMORYMAP_INFO_H__
`define __MEMORYMAP_INFO_H__


`define I_SYSTEM_SRAM_BASEADDR (32'h 40000000)
`define I_SYSTEM_SRAM_SIZE (32'h 20000)
`define I_SYSTEM_SRAM_LASTADDR (32'h 4001ffff)
`define DEFAULT_SLAVE_BASEADDR (32'h 40020000)
`define DEFAULT_SLAVE_SIZE (32'h 1000)
`define DEFAULT_SLAVE_LASTADDR (32'h 40020fff)
`define COMMON_PERI_GROUP_BASEADDR (32'h e0000000)
`define COMMON_PERI_GROUP_SIZE (32'h 10000)
`define COMMON_PERI_GROUP_LASTADDR (32'h e000ffff)
`define PLATFORM_CONTROLLER_BASEADDR (32'h e1000000)
`define PLATFORM_CONTROLLER_SIZE (32'h 40000)
`define PLATFORM_CONTROLLER_LASTADDR (32'h e103ffff)
`define EXTERNAL_PERI_GROUP_BASEADDR (32'h e1040000)
`define EXTERNAL_PERI_GROUP_SIZE (32'h 10000)
`define EXTERNAL_PERI_GROUP_LASTADDR (32'h e104ffff)
`define CORE_PERI_GROUP_BASEADDR (32'h f0000000)
`define CORE_PERI_GROUP_SIZE (32'h 1000)
`define CORE_PERI_GROUP_LASTADDR (32'h f0000fff)
`define NOC_CONTROLLER_BASEADDR (32'h 40020000)
`define IROM_BASEADDR (32'h e0000000)

`endif