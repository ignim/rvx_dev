
`define USE_SRAM
`define SRAM_HEX_SIZE 6526
`define CRM_HEX_SIZE 0
`define DRAM_HEX_SIZE 0
`define HEX_SIZE 6526