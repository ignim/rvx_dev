`ifndef __SIM_INFO_H__
`define __SIM_INFO_H__


`define SRAM_IP_INSTANCE i_system_sram
`define SRAM_WIDTH 32
`define NUM_SRAM_CELL 1
`define EXTERNAL_CLK_NAME_00 external_clk

`endif