always@(*)
begin : gen_irom_contents
rom_data = 0;
case(rom_index)
0: rom_data = 32'h e1000437;
1: rom_data = 32'h 000102b7;
2: rom_data = 32'h 02828293;
3: rom_data = 32'h 005402b3;
4: rom_data = 32'h 0002a483;
5: rom_data = 32'h e1041937;
6: rom_data = 32'h 90090913;
7: rom_data = 32'h 00010bb7;
8: rom_data = 32'h 020b8b93;
9: rom_data = 32'h 01740bb3;
10: rom_data = 32'h 000102b7;
11: rom_data = 32'h 00828293;
12: rom_data = 32'h 005402b3;
13: rom_data = 32'h 0002a303;
14: rom_data = 32'h fe030ee3;
15: rom_data = 32'h 000102b7;
16: rom_data = 32'h 005402b3;
17: rom_data = 32'h 0002a303;
18: rom_data = 32'h 00000393;
19: rom_data = 32'h 00730863;
20: rom_data = 32'h 00100393;
21: rom_data = 32'h 00730e63;
22: rom_data = 32'h 0140006f;
23: rom_data = 32'h 00200393;
24: rom_data = 32'h 000ba303;
25: rom_data = 32'h fe731ee3;
26: rom_data = 32'h 00048067;
27: rom_data = 32'h 0000006f;
28: rom_data = 32'h 000ba303;
29: rom_data = 32'h fe6014e3;
30: rom_data = 32'h 00400393;
31: rom_data = 32'h 00792023;
32: rom_data = 32'h 00300393;
33: rom_data = 32'h 00792223;
34: rom_data = 32'h 000103b7;
35: rom_data = 32'h fff38393;
36: rom_data = 32'h 00792a23;
37: rom_data = 32'h 00200393;
38: rom_data = 32'h 00792c23;
39: rom_data = 32'h 00000393;
40: rom_data = 32'h 00792823;
41: rom_data = 32'h 00100313;
42: rom_data = 32'h 00200393;
43: rom_data = 32'h 007313b3;
44: rom_data = 32'h e1041337;
45: rom_data = 32'h b5030313;
46: rom_data = 32'h 00732023;
47: rom_data = 32'h 000803b7;
48: rom_data = 32'h 04792023;
49: rom_data = 32'h 06092023;
50: rom_data = 32'h 06092223;
51: rom_data = 32'h 06092823;
52: rom_data = 32'h 00100393;
53: rom_data = 32'h 04792823;
54: rom_data = 32'h 04092a23;
55: rom_data = 32'h e10102b7;
56: rom_data = 32'h 08828293;
57: rom_data = 32'h 0002a503;
58: rom_data = 32'h 058000ef;
59: rom_data = 32'h 054000ef;
60: rom_data = 32'h 050000ef;
61: rom_data = 32'h 04c000ef;
62: rom_data = 32'h 0b4000ef;
63: rom_data = 32'h 02058e63;
64: rom_data = 32'h 00058993;
65: rom_data = 32'h 03c000ef;
66: rom_data = 32'h 038000ef;
67: rom_data = 32'h 034000ef;
68: rom_data = 32'h 030000ef;
69: rom_data = 32'h 098000ef;
70: rom_data = 32'h 00058a13;
71: rom_data = 32'h 00000593;
72: rom_data = 32'h 020000ef;
73: rom_data = 32'h 00ba0023;
74: rom_data = 32'h fff98993;
75: rom_data = 32'h 001a0a13;
76: rom_data = 32'h fe0996e3;
77: rom_data = 32'h fb5ff06f;
78: rom_data = 32'h 000ba023;
79: rom_data = 32'h f21ff06f;
80: rom_data = 32'h 00008b13;
81: rom_data = 32'h 00200393;
82: rom_data = 32'h 00792c23;
83: rom_data = 32'h 000803b7;
84: rom_data = 32'h 00838393;
85: rom_data = 32'h 04792023;
86: rom_data = 32'h 00300613;
87: rom_data = 32'h 088000ef;
88: rom_data = 32'h 01055613;
89: rom_data = 32'h 080000ef;
90: rom_data = 32'h 00855613;
91: rom_data = 32'h 078000ef;
92: rom_data = 32'h 00050613;
93: rom_data = 32'h 070000ef;
94: rom_data = 32'h 000803b7;
95: rom_data = 32'h 04792023;
96: rom_data = 32'h 064000ef;
97: rom_data = 32'h 04c92283;
98: rom_data = 32'h 01f2d313;
99: rom_data = 32'h fe031ce3;
100: rom_data = 32'h 00300393;
101: rom_data = 32'h 00792c23;
102: rom_data = 32'h 00859593;
103: rom_data = 32'h 005585b3;
104: rom_data = 32'h 00150513;
105: rom_data = 32'h 000b0093;
106: rom_data = 32'h 00008067;
107: rom_data = 32'h 0ff00293;
108: rom_data = 32'h 0055f333;
109: rom_data = 32'h 0085d593;
110: rom_data = 32'h 0055f3b3;
111: rom_data = 32'h 0085d593;
112: rom_data = 32'h 0055fe33;
113: rom_data = 32'h 0085d593;
114: rom_data = 32'h 008e1e13;
115: rom_data = 32'h 01c5e5b3;
116: rom_data = 32'h 01039393;
117: rom_data = 32'h 0075e5b3;
118: rom_data = 32'h 01831313;
119: rom_data = 32'h 0065e5b3;
120: rom_data = 32'h 00008067;
121: rom_data = 32'h 04892383;
122: rom_data = 32'h 01f3d393;
123: rom_data = 32'h fe039ce3;
124: rom_data = 32'h 04c92423;
125: rom_data = 32'h 07492383;
126: rom_data = 32'h 0013f393;
127: rom_data = 32'h fe038ce3;
128: rom_data = 32'h 00008067;
endcase
end